module main ();
    initial $display("hello, world!");
endmodule